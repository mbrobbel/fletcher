-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.UtilStr_pkg.all;
use work.UtilConv_pkg.all;

entity ProfilerStreams is
  generic (
    PROBE_COUNT_WIDTH : positive;
    OUT_COUNT_WIDTH   : positive
  );
  port (
    pcd_clk     : in  std_logic;
    pcd_reset   : in  std_logic;
    probe_valid : in  std_logic;
    probe_ready : out std_logic;
    probe_count : in  std_logic_vector(PROBE_COUNT_WIDTH-1 downto 0) := std_logic_vector(to_unsigned(1, PROBE_COUNT_WIDTH));
    enable      : in  std_logic;
    clear       : in  std_logic;
    ecount      : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    vcount      : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    rcount      : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    tcount      : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0);
    pcount      : out std_logic_vector(OUT_COUNT_WIDTH-1 downto 0)
  );
end ProfilerStreams;

architecture Behavioral of ProfilerStreams is
begin

  t_count_proc: process is
    variable transfers : natural := 0;
  begin
    -- Wait for reset.
    loop
      wait until rising_edge(pcd_clk) ;
      exit when pcd_reset = '0';
    end loop;
    
    if (enable = '1') then
      loop
        wait until rising_edge(pcd_clk);
        exit when probe_valid = '1' and probe_ready = '1';
      end loop;
      
      transfers := transfers + 1;
      
      tcount <= std_logic_vector(to_unsigned(transfers, 32));    
      
      println("Transfers: " & slvToDec(tcount));
    end if;
  end process;

end architecture;
